library verilog;
use verilog.vl_types.all;
entity mp3_top_sv_unit is
end mp3_top_sv_unit;
