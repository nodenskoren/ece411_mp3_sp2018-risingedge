library verilog;
use verilog.vl_types.all;
library work;
entity EX_MEM_pipeline is
    port(
        clk             : in     vl_logic;
        is_j_in         : in     vl_logic;
        alu_out_in      : in     vl_logic_vector(15 downto 0);
        addr_adder_out_in: in     vl_logic_vector(15 downto 0);
        pc_in           : in     vl_logic_vector(15 downto 0);
        dest_in         : in     vl_logic_vector(2 downto 0);
        nzp_in          : in     vl_logic_vector(2 downto 0);
        is_br_in        : in     vl_logic;
        is_jsr_in       : in     vl_logic;
        is_trap_in      : in     vl_logic;
        load_cc_in      : in     vl_logic;
        load_regfile_in : in     vl_logic;
        mem_read_in     : in     vl_logic;
        mem_write_in    : in     vl_logic;
        regfilemux_sel_in: in     vl_logic_vector(2 downto 0);
        dest_data_in    : in     vl_logic_vector(15 downto 0);
        trapvector_in   : in     vl_logic_vector(15 downto 0);
        addr_sel_in     : in     vl_logic_vector(1 downto 0);
        mem_byte_enable_in: in     vl_logic_vector(1 downto 0);
        is_ldi_in       : in     vl_logic;
        is_sti_in       : in     vl_logic;
        ctrl_in         : in     work.lc3b_types.lc3b_control_word;
        is_ldb_stb_in   : in     vl_logic;
        is_j_out        : out    vl_logic;
        alu_out_out     : out    vl_logic_vector(15 downto 0);
        addr_adder_out_out: out    vl_logic_vector(15 downto 0);
        pc_out          : out    vl_logic_vector(15 downto 0);
        dest_out        : out    vl_logic_vector(2 downto 0);
        nzp_out         : out    vl_logic_vector(2 downto 0);
        is_br_out       : out    vl_logic;
        load_cc_out     : out    vl_logic;
        load_regfile_out: out    vl_logic;
        mem_read_out    : out    vl_logic;
        mem_write_out   : out    vl_logic;
        regfilemux_sel_out: out    vl_logic_vector(2 downto 0);
        dest_data_out   : out    vl_logic_vector(15 downto 0);
        is_jsr_out      : out    vl_logic;
        is_trap_out     : out    vl_logic;
        trapvector_out  : out    vl_logic_vector(15 downto 0);
        addr_sel_out    : out    vl_logic_vector(1 downto 0);
        mem_byte_enable_out: out    vl_logic_vector(1 downto 0);
        is_ldi_out      : out    vl_logic;
        is_sti_out      : out    vl_logic;
        ctrl_out        : out    work.lc3b_types.lc3b_control_word;
        is_ldb_stb_out  : out    vl_logic;
        operation_in    : in     work.lc3b_types.lc3b_opcode;
        operation_out   : out    work.lc3b_types.lc3b_opcode;
        instruction_in  : in     vl_logic_vector(15 downto 0);
        instruction_out : out    vl_logic_vector(15 downto 0);
        stall_pipeline  : in     vl_logic;
        branch_history_in: in     vl_logic_vector(7 downto 0);
        branch_history_out: out    vl_logic_vector(7 downto 0);
        branch_prediction_in: in     vl_logic;
        branch_prediction_out: out    vl_logic;
        branch_address_in: in     vl_logic_vector(15 downto 0);
        branch_address_out: out    vl_logic_vector(15 downto 0)
    );
end EX_MEM_pipeline;
