library verilog;
use verilog.vl_types.all;
entity forwarding_unit_2_sv_unit is
end forwarding_unit_2_sv_unit;
