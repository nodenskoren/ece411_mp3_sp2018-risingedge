library verilog;
use verilog.vl_types.all;
entity cache_prefetch_sv_unit is
end cache_prefetch_sv_unit;
