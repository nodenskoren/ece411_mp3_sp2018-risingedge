library verilog;
use verilog.vl_types.all;
entity counter_decoder_sv_unit is
end counter_decoder_sv_unit;
