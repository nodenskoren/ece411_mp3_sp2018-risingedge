library verilog;
use verilog.vl_types.all;
entity set_sel_sv_unit is
end set_sel_sv_unit;
