library verilog;
use verilog.vl_types.all;
entity EX_MEM_pipeline_sv_unit is
end EX_MEM_pipeline_sv_unit;
