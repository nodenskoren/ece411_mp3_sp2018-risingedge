library verilog;
use verilog.vl_types.all;
entity stall_unit_2_sv_unit is
end stall_unit_2_sv_unit;
