library verilog;
use verilog.vl_types.all;
entity mp3_top is
end mp3_top;
