library verilog;
use verilog.vl_types.all;
entity cache_control4way_sv_unit is
end cache_control4way_sv_unit;
