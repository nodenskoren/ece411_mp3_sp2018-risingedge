library verilog;
use verilog.vl_types.all;
entity cache_datapath_prefetch_sv_unit is
end cache_datapath_prefetch_sv_unit;
