library verilog;
use verilog.vl_types.all;
entity stall_unit_sv_unit is
end stall_unit_sv_unit;
