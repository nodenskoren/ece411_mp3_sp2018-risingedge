library verilog;
use verilog.vl_types.all;
entity magic_memory is
end magic_memory;
