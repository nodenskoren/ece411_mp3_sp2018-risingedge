library verilog;
use verilog.vl_types.all;
entity l2cache is
end l2cache;
