library verilog;
use verilog.vl_types.all;
entity zextadj_sv_unit is
end zextadj_sv_unit;
