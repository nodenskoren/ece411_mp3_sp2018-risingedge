library verilog;
use verilog.vl_types.all;
entity evict_buffer_sv_unit is
end evict_buffer_sv_unit;
