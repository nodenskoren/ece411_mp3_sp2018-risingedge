library verilog;
use verilog.vl_types.all;
entity always_branch_sv_unit is
end always_branch_sv_unit;
