library verilog;
use verilog.vl_types.all;
entity wb_interconnect_sv_unit is
end wb_interconnect_sv_unit;
