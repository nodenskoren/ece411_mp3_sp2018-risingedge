library verilog;
use verilog.vl_types.all;
entity l1arbiter_sv_unit is
end l1arbiter_sv_unit;
