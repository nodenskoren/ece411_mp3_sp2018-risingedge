library verilog;
use verilog.vl_types.all;
entity cache_control_prefetch_sv_unit is
end cache_control_prefetch_sv_unit;
