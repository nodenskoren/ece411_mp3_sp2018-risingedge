library verilog;
use verilog.vl_types.all;
entity cache_writeword_sv_unit is
end cache_writeword_sv_unit;
