library verilog;
use verilog.vl_types.all;
entity zext4_sv_unit is
end zext4_sv_unit;
