library verilog;
use verilog.vl_types.all;
entity pseudoLRU4way_sv_unit is
end pseudoLRU4way_sv_unit;
