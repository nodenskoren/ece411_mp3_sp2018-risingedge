library verilog;
use verilog.vl_types.all;
entity line_to_word_sv_unit is
end line_to_word_sv_unit;
