library verilog;
use verilog.vl_types.all;
entity wb_interconnect is
end wb_interconnect;
