library verilog;
use verilog.vl_types.all;
entity branch_unit_sv_unit is
end branch_unit_sv_unit;
