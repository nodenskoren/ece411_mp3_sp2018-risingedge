library verilog;
use verilog.vl_types.all;
entity sext5_sv_unit is
end sext5_sv_unit;
