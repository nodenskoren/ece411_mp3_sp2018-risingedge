library verilog;
use verilog.vl_types.all;
entity l2cache4way_sv_unit is
end l2cache4way_sv_unit;
