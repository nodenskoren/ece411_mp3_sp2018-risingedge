library verilog;
use verilog.vl_types.all;
entity wishbone is
    port(
        CLK             : in     vl_logic
    );
end wishbone;
