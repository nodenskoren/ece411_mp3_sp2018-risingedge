library verilog;
use verilog.vl_types.all;
entity static_branch_prediction_sv_unit is
end static_branch_prediction_sv_unit;
