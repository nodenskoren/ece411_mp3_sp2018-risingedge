library verilog;
use verilog.vl_types.all;
entity l2cache_sv_unit is
end l2cache_sv_unit;
