library verilog;
use verilog.vl_types.all;
entity counter_control_sv_unit is
end counter_control_sv_unit;
