library verilog;
use verilog.vl_types.all;
entity cache_datapath4way_sv_unit is
end cache_datapath4way_sv_unit;
